----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    19:48:40 11/30/2017 
-- Design Name: 
-- Module Name:    DecROB - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity DecROB is
Port ( InD : in  STD_LOGIC_VECTOR (2 downto 0);
           OutD : out  STD_LOGIC_VECTOR (7 downto 0));
end DecROB;

architecture Behavioral of DecROB is

begin


with InD select
			OutD <= "00000000" when "000",--EDW KAI TO KOLPO TOU R0=0
					  "00000010" when "001",
					  "00000100" when "010",
					  "00001000" when "011",
					  "00010000" when "100",
					  "00100000" when "101",
					  "01000000" when "110",
					  "10000000" when others;
					 

end Behavioral;

